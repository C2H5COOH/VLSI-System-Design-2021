// `include "../AXI/AXI_slave/AXISlave.sv"
`include "AXI/AXI_slave_SRAM/AXISlaveSRAM.sv"

module SRAM_wrapper (
  input clock,
	input reset,
  // READ ADDRESS
	input [`AXI_IDS_BITS-1:0] ARID,
	input [`AXI_ADDR_BITS-1:0] ARADDR,
	input [`AXI_LEN_BITS-1:0] ARLEN,
	input [`AXI_SIZE_BITS-1:0] ARSIZE,
	input [`AXI_BURST_BITS-1:0] ARBURST,
	input ARVALID,
	output ARREADY,
	// READ DATA
	output [`AXI_IDS_BITS-1:0] RID,
	output [`AXI_DATA_BITS-1:0] RDATA,
	output [`AXI_RESP_BITS-1:0] RRESP,
	output RLAST,
	output RVALID,
	input RREADY,
    // WRITE ADDRESS
	input [`AXI_IDS_BITS-1:0] AWID,
	input [`AXI_ADDR_BITS-1:0] AWADDR,
	input [`AXI_LEN_BITS-1:0] AWLEN,
	input [`AXI_SIZE_BITS-1:0] AWSIZE,
	input [`AXI_BURST_BITS-1:0] AWBURST,
	input AWVALID,
	output AWREADY,
	// WRITE DATA
	input [`AXI_DATA_BITS-1:0] WDATA,
	input [`AXI_STRB_BITS-1:0] WSTRB,
	input WLAST,
	input WVALID,
	output WREADY,
	// WRITE RESPONSE
	output [`AXI_IDS_BITS-1:0] BID,
	output [`AXI_RESP_BITS-1:0] BRESP,
	output BVALID,
	input BREADY
);
  // Wire
  logic [`AXI_ADDR_BITS-1:0] Address;
  logic CS;
  logic OE;
  logic [`AXI_STRB_BITS-1:0] WEB;
  logic [12:0] A;
  logic [`AXI_DATA_BITS-1:0] DI;
  logic [`AXI_DATA_BITS-1:0] DO;

  // Module
  AXISlaveSRAM axiSlaveSRAM
  (
    .clock(clock),
    .reset(reset),
      // READ ADDRESS
    .ARID(ARID),
    .ARADDR(ARADDR),
    .ARLEN(ARLEN),
    .ARSIZE(ARSIZE),
    .ARBURST(ARBURST),
    .ARVALID(ARVALID),
    .ARREADY(ARREADY),
    // READ DATA
    .RID(RID),
    .RDATA(RDATA),
    .RRESP(RRESP),
    .RLAST(RLAST),
    .RVALID(RVALID),
    .RREADY(RREADY),
      // WRITE ADDRESS
    .AWID(AWID),
    .AWADDR(AWADDR),
    .AWLEN(AWLEN),
    .AWSIZE(AWSIZE),
    .AWBURST(AWBURST),
    .AWVALID(AWVALID),
    .AWREADY(AWREADY),
    // WRITE DATA
    .WDATA(WDATA),
    .WSTRB(WSTRB),
    .WLAST(WLAST),
    .WVALID(WVALID),
    .WREADY(WREADY),
    // WRITE RESPONSE
    .BID(BID),
    .BRESP(BRESP),
    .BVALID(BVALID),
    .BREADY(BREADY),
    // Slave
    .Address(Address),
    .ReadEnable(OE),
    .DataRead(DO),
    .WriteEnable(WEB),
    .DataWrite(DI)
  );
  SRAM_64 i_SRAM 
  (
    .A0   (A[0]  ),
    .A1   (A[1]  ),
    .A2   (A[2]  ),
    .A3   (A[3]  ),
    .A4   (A[4]  ),
    .A5   (A[5]  ),
    .A6   (A[6]  ),
    .A7   (A[7]  ),
    .A8   (A[8]  ),
    .A9   (A[9]  ),
    .A10  (A[10] ),
    .A11  (A[11] ),
    .A12  (A[12] ),

    .DO0  (DO[0] ),
    .DO1  (DO[1] ),
    .DO2  (DO[2] ),
    .DO3  (DO[3] ),
    .DO4  (DO[4] ),
    .DO5  (DO[5] ),
    .DO6  (DO[6] ),
    .DO7  (DO[7] ),
    .DO8  (DO[8] ),
    .DO9  (DO[9] ),
    .DO10 (DO[10]),
    .DO11 (DO[11]),
    .DO12 (DO[12]),
    .DO13 (DO[13]),
    .DO14 (DO[14]),
    .DO15 (DO[15]),
    .DO16 (DO[16]),
    .DO17 (DO[17]),
    .DO18 (DO[18]),
    .DO19 (DO[19]),
    .DO20 (DO[20]),
    .DO21 (DO[21]),
    .DO22 (DO[22]),
    .DO23 (DO[23]),
    .DO24 (DO[24]),
    .DO25 (DO[25]),
    .DO26 (DO[26]),
    .DO27 (DO[27]),
    .DO28 (DO[28]),
    .DO29 (DO[29]),
    .DO30 (DO[30]),
    .DO31 (DO[31]),
    .DO32 (DO[32]),
    .DO33 (DO[33]),
    .DO34 (DO[34]),
    .DO35 (DO[35]),
    .DO36 (DO[36]),
    .DO37 (DO[37]),
    .DO38 (DO[38]),
    .DO39 (DO[39]),
    .DO40 (DO[40]),
    .DO41 (DO[41]),
    .DO42 (DO[42]),
    .DO43 (DO[43]),
    .DO44 (DO[44]),
    .DO45 (DO[45]),
    .DO46 (DO[46]),
    .DO47 (DO[47]),
    .DO48 (DO[48]),
    .DO49 (DO[49]),
    .DO50 (DO[50]),
    .DO51 (DO[51]),
    .DO52 (DO[52]),
    .DO53 (DO[53]),
    .DO54 (DO[54]),
    .DO55 (DO[55]),
    .DO56 (DO[56]),
    .DO57 (DO[57]),
    .DO58 (DO[58]),
    .DO59 (DO[59]),
    .DO60 (DO[60]),
    .DO61 (DO[61]),
    .DO62 (DO[62]),
    .DO63 (DO[63]),
    .DI0  (DI[0] ),
    .DI1  (DI[1] ),
    .DI2  (DI[2] ),
    .DI3  (DI[3] ),
    .DI4  (DI[4] ),
    .DI5  (DI[5] ),
    .DI6  (DI[6] ),
    .DI7  (DI[7] ),
    .DI8  (DI[8] ),
    .DI9  (DI[9] ),
    .DI10 (DI[10]),
    .DI11 (DI[11]),
    .DI12 (DI[12]),
    .DI13 (DI[13]),
    .DI14 (DI[14]),
    .DI15 (DI[15]),
    .DI16 (DI[16]),
    .DI17 (DI[17]),
    .DI18 (DI[18]),
    .DI19 (DI[19]),
    .DI20 (DI[20]),
    .DI21 (DI[21]),
    .DI22 (DI[22]),
    .DI23 (DI[23]),
    .DI24 (DI[24]),
    .DI25 (DI[25]),
    .DI26 (DI[26]),
    .DI27 (DI[27]),
    .DI28 (DI[28]),
    .DI29 (DI[29]),
    .DI30 (DI[30]),
    .DI31 (DI[31]),
    .DI32 (DI[32]),
    .DI33 (DI[33]),
    .DI34 (DI[34]),
    .DI35 (DI[35]),
    .DI36 (DI[36]),
    .DI37 (DI[37]),
    .DI38 (DI[38]),
    .DI39 (DI[39]),
    .DI40 (DI[40]),
    .DI41 (DI[41]),
    .DI42 (DI[42]),
    .DI43 (DI[43]),
    .DI44 (DI[44]),
    .DI45 (DI[45]),
    .DI46 (DI[46]),
    .DI47 (DI[47]),
    .DI48 (DI[48]),
    .DI49 (DI[49]),
    .DI50 (DI[50]),
    .DI51 (DI[51]),
    .DI52 (DI[52]),
    .DI53 (DI[53]),
    .DI54 (DI[54]),
    .DI55 (DI[55]),
    .DI56 (DI[56]),
    .DI57 (DI[57]),
    .DI58 (DI[58]),
    .DI59 (DI[59]),
    .DI60 (DI[60]),
    .DI61 (DI[61]),
    .DI62 (DI[62]),
    .DI63 (DI[63]),
    .CK   (clock),
    .WEB0 (WEB[0]),
    .WEB1 (WEB[1]),
    .WEB2 (WEB[2]),
    .WEB3 (WEB[3]),
    .WEB4 (WEB[4]),
    .WEB5 (WEB[5]),
    .WEB6 (WEB[6]),
    .WEB7 (WEB[7]),
    .OE   (OE    ),
    .CS   (CS    )
  );

  assign A = Address[15:3];
  assign CS = 1'b1;
endmodule
