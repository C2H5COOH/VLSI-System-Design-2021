`ifndef CONFIG_SVH
`define CONFIG_SVH

`define DATA_BIT_WIDTH 32
`define REGISTER_NUM   32

`endif

