`include "TPU_def.svh"

module OFM_wrapper (
    input                           CK,
    input [`OFM_SRAM_ADDR_BIT-1:0]  A,
    input [`MAC_OUT_BIT-1:0]        DI  [0:`SYS_WIDTH-1],
    input [`SYS_WIDTH-1:0]          WEB,
    input                           OE,
    input                           CS,
    output logic [`MAC_OUT_BIT-1:0] DO  [0:`SYS_WIDTH-1]
);
SUMA180_464X24X4BM1 iSRAM24x4_0 (
    .A0(A[0]),
    .A1(A[1]),
    .A2(A[2]),
    .A3(A[3]),
    .A4(A[4]),
    .A5(A[5]),
    .A6(A[6]),
    .A7(A[7]),
    .A8(A[8]),
    .DO0 (DO[0][0]),
    .DO1 (DO[0][1]),
    .DO2 (DO[0][2]),
    .DO3 (DO[0][3]),
    .DO4 (DO[0][4]),
    .DO5 (DO[0][5]),
    .DO6 (DO[0][6]),
    .DO7 (DO[0][7]),
    .DO8 (DO[0][8]),
    .DO9 (DO[0][9]),
    .DO10(DO[0][10]),
    .DO11(DO[0][11]),
    .DO12(DO[0][12]),
    .DO13(DO[0][13]),
    .DO14(DO[0][14]),
    .DO15(DO[0][15]),
    .DO16(DO[0][16]),
    .DO17(DO[0][17]),
    .DO18(DO[0][18]),
    .DO19(DO[0][19]),
    .DO20(DO[0][20]),
    .DO21(DO[0][21]),
    .DO22(DO[0][22]),
    .DO23(DO[0][23]),
    .DO24(DO[1][0]),
    .DO25(DO[1][1]),
    .DO26(DO[1][2]),
    .DO27(DO[1][3]),
    .DO28(DO[1][4]),
    .DO29(DO[1][5]),
    .DO30(DO[1][6]),
    .DO31(DO[1][7]),
    .DO32(DO[1][8]),
    .DO33(DO[1][9]),
    .DO34(DO[1][10]),
    .DO35(DO[1][11]),
    .DO36(DO[1][12]),
    .DO37(DO[1][13]),
    .DO38(DO[1][14]),
    .DO39(DO[1][15]),
    .DO40(DO[1][16]),
    .DO41(DO[1][17]),
    .DO42(DO[1][18]),
    .DO43(DO[1][19]),
    .DO44(DO[1][20]),
    .DO45(DO[1][21]),
    .DO46(DO[1][22]),
    .DO47(DO[1][23]),
    .DO48(DO[2][0]),
    .DO49(DO[2][1]),
    .DO50(DO[2][2]),
    .DO51(DO[2][3]),
    .DO52(DO[2][4]),
    .DO53(DO[2][5]),
    .DO54(DO[2][6]),
    .DO55(DO[2][7]),
    .DO56(DO[2][8]),
    .DO57(DO[2][9]),
    .DO58(DO[2][10]),
    .DO59(DO[2][11]),
    .DO60(DO[2][12]),
    .DO61(DO[2][13]),
    .DO62(DO[2][14]),
    .DO63(DO[2][15]),
    .DO64(DO[2][16]),
    .DO65(DO[2][17]),
    .DO66(DO[2][18]),
    .DO67(DO[2][19]),
    .DO68(DO[2][20]),
    .DO69(DO[2][21]),
    .DO70(DO[2][22]),
    .DO71(DO[2][23]),
    .DO72(DO[3][0]),
    .DO73(DO[3][1]),
    .DO74(DO[3][2]),
    .DO75(DO[3][3]),
    .DO76(DO[3][4]),
    .DO77(DO[3][5]),
    .DO78(DO[3][6]),
    .DO79(DO[3][7]),
    .DO80(DO[3][8]),
    .DO81(DO[3][9]),
    .DO82(DO[3][10]),
    .DO83(DO[3][11]),
    .DO84(DO[3][12]),
    .DO85(DO[3][13]),
    .DO86(DO[3][14]),
    .DO87(DO[3][15]),
    .DO88(DO[3][16]),
    .DO89(DO[3][17]),
    .DO90(DO[3][18]),
    .DO91(DO[3][19]),
    .DO92(DO[3][20]),
    .DO93(DO[3][21]),
    .DO94(DO[3][22]),
    .DO95(DO[3][23]),
    .DI0 (DI[0][0]),
    .DI1 (DI[0][1]),
    .DI2 (DI[0][2]),
    .DI3 (DI[0][3]),
    .DI4 (DI[0][4]),
    .DI5 (DI[0][5]),
    .DI6 (DI[0][6]),
    .DI7 (DI[0][7]),
    .DI8 (DI[0][8]),
    .DI9 (DI[0][9]),
    .DI10(DI[0][10]),
    .DI11(DI[0][11]),
    .DI12(DI[0][12]),
    .DI13(DI[0][13]),
    .DI14(DI[0][14]),
    .DI15(DI[0][15]),
    .DI16(DI[0][16]),
    .DI17(DI[0][17]),
    .DI18(DI[0][18]),
    .DI19(DI[0][19]),
    .DI20(DI[0][20]),
    .DI21(DI[0][21]),
    .DI22(DI[0][22]),
    .DI23(DI[0][23]),
    .DI24(DI[1][0]),
    .DI25(DI[1][1]),
    .DI26(DI[1][2]),
    .DI27(DI[1][3]),
    .DI28(DI[1][4]),
    .DI29(DI[1][5]),
    .DI30(DI[1][6]),
    .DI31(DI[1][7]),
    .DI32(DI[1][8]),
    .DI33(DI[1][9]),
    .DI34(DI[1][10]),
    .DI35(DI[1][11]),
    .DI36(DI[1][12]),
    .DI37(DI[1][13]),
    .DI38(DI[1][14]),
    .DI39(DI[1][15]),
    .DI40(DI[1][16]),
    .DI41(DI[1][17]),
    .DI42(DI[1][18]),
    .DI43(DI[1][19]),
    .DI44(DI[1][20]),
    .DI45(DI[1][21]),
    .DI46(DI[1][22]),
    .DI47(DI[1][23]),
    .DI48(DI[2][0]),
    .DI49(DI[2][1]),
    .DI50(DI[2][2]),
    .DI51(DI[2][3]),
    .DI52(DI[2][4]),
    .DI53(DI[2][5]),
    .DI54(DI[2][6]),
    .DI55(DI[2][7]),
    .DI56(DI[2][8]),
    .DI57(DI[2][9]),
    .DI58(DI[2][10]),
    .DI59(DI[2][11]),
    .DI60(DI[2][12]),
    .DI61(DI[2][13]),
    .DI62(DI[2][14]),
    .DI63(DI[2][15]),
    .DI64(DI[2][16]),
    .DI65(DI[2][17]),
    .DI66(DI[2][18]),
    .DI67(DI[2][19]),
    .DI68(DI[2][20]),
    .DI69(DI[2][21]),
    .DI70(DI[2][22]),
    .DI71(DI[2][23]),
    .DI72(DI[3][0]),
    .DI73(DI[3][1]),
    .DI74(DI[3][2]),
    .DI75(DI[3][3]),
    .DI76(DI[3][4]),
    .DI77(DI[3][5]),
    .DI78(DI[3][6]),
    .DI79(DI[3][7]),
    .DI80(DI[3][8]),
    .DI81(DI[3][9]),
    .DI82(DI[3][10]),
    .DI83(DI[3][11]),
    .DI84(DI[3][12]),
    .DI85(DI[3][13]),
    .DI86(DI[3][14]),
    .DI87(DI[3][15]),
    .DI88(DI[3][16]),
    .DI89(DI[3][17]),
    .DI90(DI[3][18]),
    .DI91(DI[3][19]),
    .DI92(DI[3][20]),
    .DI93(DI[3][21]),
    .DI94(DI[3][22]),
    .DI95(DI[3][23]),
    .CK(CK),
    .WEB0(WEB[0]),
    .WEB1(WEB[1]),
    .WEB2(WEB[2]),
    .WEB3(WEB[3]),
    .OE(OE),
    .CS(CS)
);

SUMA180_464X24X4BM1 iSRAM24x4_1 (
    .A0(A[0]),
    .A1(A[1]),
    .A2(A[2]),
    .A3(A[3]),
    .A4(A[4]),
    .A5(A[5]),
    .A6(A[6]),
    .A7(A[7]),
    .A8(A[8]),
    .DO0 (DO[4][0]),
    .DO1 (DO[4][1]),
    .DO2 (DO[4][2]),
    .DO3 (DO[4][3]),
    .DO4 (DO[4][4]),
    .DO5 (DO[4][5]),
    .DO6 (DO[4][6]),
    .DO7 (DO[4][7]),
    .DO8 (DO[4][8]),
    .DO9 (DO[4][9]),
    .DO10(DO[4][10]),
    .DO11(DO[4][11]),
    .DO12(DO[4][12]),
    .DO13(DO[4][13]),
    .DO14(DO[4][14]),
    .DO15(DO[4][15]),
    .DO16(DO[4][16]),
    .DO17(DO[4][17]),
    .DO18(DO[4][18]),
    .DO19(DO[4][19]),
    .DO20(DO[4][20]),
    .DO21(DO[4][21]),
    .DO22(DO[4][22]),
    .DO23(DO[4][23]),
    .DO24(DO[5][0]),
    .DO25(DO[5][1]),
    .DO26(DO[5][2]),
    .DO27(DO[5][3]),
    .DO28(DO[5][4]),
    .DO29(DO[5][5]),
    .DO30(DO[5][6]),
    .DO31(DO[5][7]),
    .DO32(DO[5][8]),
    .DO33(DO[5][9]),
    .DO34(DO[5][10]),
    .DO35(DO[5][11]),
    .DO36(DO[5][12]),
    .DO37(DO[5][13]),
    .DO38(DO[5][14]),
    .DO39(DO[5][15]),
    .DO40(DO[5][16]),
    .DO41(DO[5][17]),
    .DO42(DO[5][18]),
    .DO43(DO[5][19]),
    .DO44(DO[5][20]),
    .DO45(DO[5][21]),
    .DO46(DO[5][22]),
    .DO47(DO[5][23]),
    .DO48(DO[6][0]),
    .DO49(DO[6][1]),
    .DO50(DO[6][2]),
    .DO51(DO[6][3]),
    .DO52(DO[6][4]),
    .DO53(DO[6][5]),
    .DO54(DO[6][6]),
    .DO55(DO[6][7]),
    .DO56(DO[6][8]),
    .DO57(DO[6][9]),
    .DO58(DO[6][10]),
    .DO59(DO[6][11]),
    .DO60(DO[6][12]),
    .DO61(DO[6][13]),
    .DO62(DO[6][14]),
    .DO63(DO[6][15]),
    .DO64(DO[6][16]),
    .DO65(DO[6][17]),
    .DO66(DO[6][18]),
    .DO67(DO[6][19]),
    .DO68(DO[6][20]),
    .DO69(DO[6][21]),
    .DO70(DO[6][22]),
    .DO71(DO[6][23]),
    .DO72(DO[7][0]),
    .DO73(DO[7][1]),
    .DO74(DO[7][2]),
    .DO75(DO[7][3]),
    .DO76(DO[7][4]),
    .DO77(DO[7][5]),
    .DO78(DO[7][6]),
    .DO79(DO[7][7]),
    .DO80(DO[7][8]),
    .DO81(DO[7][9]),
    .DO82(DO[7][10]),
    .DO83(DO[7][11]),
    .DO84(DO[7][12]),
    .DO85(DO[7][13]),
    .DO86(DO[7][14]),
    .DO87(DO[7][15]),
    .DO88(DO[7][16]),
    .DO89(DO[7][17]),
    .DO90(DO[7][18]),
    .DO91(DO[7][19]),
    .DO92(DO[7][20]),
    .DO93(DO[7][21]),
    .DO94(DO[7][22]),
    .DO95(DO[7][23]),
    .DI0 (DI[4][0]),
    .DI1 (DI[4][1]),
    .DI2 (DI[4][2]),
    .DI3 (DI[4][3]),
    .DI4 (DI[4][4]),
    .DI5 (DI[4][5]),
    .DI6 (DI[4][6]),
    .DI7 (DI[4][7]),
    .DI8 (DI[4][8]),
    .DI9 (DI[4][9]),
    .DI10(DI[4][10]),
    .DI11(DI[4][11]),
    .DI12(DI[4][12]),
    .DI13(DI[4][13]),
    .DI14(DI[4][14]),
    .DI15(DI[4][15]),
    .DI16(DI[4][16]),
    .DI17(DI[4][17]),
    .DI18(DI[4][18]),
    .DI19(DI[4][19]),
    .DI20(DI[4][20]),
    .DI21(DI[4][21]),
    .DI22(DI[4][22]),
    .DI23(DI[4][23]),
    .DI24(DI[5][0]),
    .DI25(DI[5][1]),
    .DI26(DI[5][2]),
    .DI27(DI[5][3]),
    .DI28(DI[5][4]),
    .DI29(DI[5][5]),
    .DI30(DI[5][6]),
    .DI31(DI[5][7]),
    .DI32(DI[5][8]),
    .DI33(DI[5][9]),
    .DI34(DI[5][10]),
    .DI35(DI[5][11]),
    .DI36(DI[5][12]),
    .DI37(DI[5][13]),
    .DI38(DI[5][14]),
    .DI39(DI[5][15]),
    .DI40(DI[5][16]),
    .DI41(DI[5][17]),
    .DI42(DI[5][18]),
    .DI43(DI[5][19]),
    .DI44(DI[5][20]),
    .DI45(DI[5][21]),
    .DI46(DI[5][22]),
    .DI47(DI[5][23]),
    .DI48(DI[6][0]),
    .DI49(DI[6][1]),
    .DI50(DI[6][2]),
    .DI51(DI[6][3]),
    .DI52(DI[6][4]),
    .DI53(DI[6][5]),
    .DI54(DI[6][6]),
    .DI55(DI[6][7]),
    .DI56(DI[6][8]),
    .DI57(DI[6][9]),
    .DI58(DI[6][10]),
    .DI59(DI[6][11]),
    .DI60(DI[6][12]),
    .DI61(DI[6][13]),
    .DI62(DI[6][14]),
    .DI63(DI[6][15]),
    .DI64(DI[6][16]),
    .DI65(DI[6][17]),
    .DI66(DI[6][18]),
    .DI67(DI[6][19]),
    .DI68(DI[6][20]),
    .DI69(DI[6][21]),
    .DI70(DI[6][22]),
    .DI71(DI[6][23]),
    .DI72(DI[7][0]),
    .DI73(DI[7][1]),
    .DI74(DI[7][2]),
    .DI75(DI[7][3]),
    .DI76(DI[7][4]),
    .DI77(DI[7][5]),
    .DI78(DI[7][6]),
    .DI79(DI[7][7]),
    .DI80(DI[7][8]),
    .DI81(DI[7][9]),
    .DI82(DI[7][10]),
    .DI83(DI[7][11]),
    .DI84(DI[7][12]),
    .DI85(DI[7][13]),
    .DI86(DI[7][14]),
    .DI87(DI[7][15]),
    .DI88(DI[7][16]),
    .DI89(DI[7][17]),
    .DI90(DI[7][18]),
    .DI91(DI[7][19]),
    .DI92(DI[7][20]),
    .DI93(DI[7][21]),
    .DI94(DI[7][22]),
    .DI95(DI[7][23]),
    .CK(CK),
    .WEB0(WEB[4]),
    .WEB1(WEB[5]),
    .WEB2(WEB[6]),
    .WEB3(WEB[7]),
    .OE(OE),
    .CS(CS)
);
endmodule