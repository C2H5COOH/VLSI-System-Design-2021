//================================================
// Auther:      Chang Wan-Yun (Claire)
// Filename:    AXI.sv
// Description: Top module of AXI
// Version:     1.0 
//================================================
`include "AXI_def.svh"
`include "AXI_rd.sv"
`include "AXI_wr.sv"

module AXI(
    input ACLK,
    input ARESETn,
    //MASTER INTERFACE
    // M0
    // READ
    input [`AXI_ID_BITS-1:0]          ARID_M0,
    input [`AXI_ADDR_BITS-1:0]        ARADDR_M0,
    input [`AXI_LEN_BITS-1:0]         ARLEN_M0,
    input [`AXI_SIZE_BITS-1:0]        ARSIZE_M0,
    input [`AXI_BURST_BITS-1:0]       ARBURST_M0,
    input                             ARVALID_M0,
    output logic                      ARREADY_M0,
    output logic [`AXI_ID_BITS-1:0]   RID_M0,
    output logic [`AXI_DATA_BITS-1:0] RDATA_M0,
    output logic [`AXI_RESP_BITS-1:0] RRESP_M0,
    output logic                      RLAST_M0,
    output logic                      RVALID_M0,
    input                             RREADY_M0,
    // M1
    // WRITE
    input [`AXI_ID_BITS-1:0]          AWID_M1,
    input [`AXI_ADDR_BITS-1:0]        AWADDR_M1,
    input [`AXI_LEN_BITS-1:0]         AWLEN_M1,
    input [`AXI_SIZE_BITS-1:0]        AWSIZE_M1,
    input [`AXI_BURST_BITS-1:0]       AWBURST_M1,
    input                             AWVALID_M1,
    output logic                      AWREADY_M1,
    input [`AXI_DATA_BITS-1:0]        WDATA_M1,
    input [`AXI_STRB_BITS-1:0]        WSTRB_M1,
    input                             WLAST_M1,
    input                             WVALID_M1,
    output logic                      WREADY_M1,
    output logic [`AXI_ID_BITS-1:0]   BID_M1,
    output logic [`AXI_RESP_BITS-1:0] BRESP_M1,
    output logic                      BVALID_M1,
    input                             BREADY_M1,
    // READ
    input [`AXI_ID_BITS-1:0]          ARID_M1,
    input [`AXI_ADDR_BITS-1:0]        ARADDR_M1,
    input [`AXI_LEN_BITS-1:0]         ARLEN_M1,
    input [`AXI_SIZE_BITS-1:0]        ARSIZE_M1,
    input [`AXI_BURST_BITS-1:0]       ARBURST_M1,
    input                             ARVALID_M1,
    output logic                      ARREADY_M1,
    output logic [`AXI_ID_BITS-1:0]   RID_M1,
    output logic [`AXI_DATA_BITS-1:0] RDATA_M1,
    output logic [`AXI_RESP_BITS-1:0] RRESP_M1,
    output logic                      RLAST_M1,
    output logic                      RVALID_M1,
    input                             RREADY_M1,
    // M2
    // WRITE
    input [`AXI_ID_BITS-1:0]          AWID_M2,
    input [`AXI_ADDR_BITS-1:0]        AWADDR_M2,
    input [`AXI_LEN_BITS-1:0]         AWLEN_M2,
    input [`AXI_SIZE_BITS-1:0]        AWSIZE_M2,
    input [`AXI_BURST_BITS-1:0]       AWBURST_M2,
    input                             AWVALID_M2,
    output logic                      AWREADY_M2,
    input [`AXI_DATA_BITS-1:0]        WDATA_M2,
    input [`AXI_STRB_BITS-1:0]        WSTRB_M2,
    input                             WLAST_M2,
    input                             WVALID_M2,
    output logic                      WREADY_M2,
    output logic [`AXI_ID_BITS-1:0]   BID_M2,
    output logic [`AXI_RESP_BITS-1:0] BRESP_M2,
    output logic                      BVALID_M2,
    input                             BREADY_M2,
    // READ
    input [`AXI_ID_BITS-1:0]          ARID_M2,
    input [`AXI_ADDR_BITS-1:0]        ARADDR_M2,
    input [`AXI_LEN_BITS-1:0]         ARLEN_M2,
    input [`AXI_SIZE_BITS-1:0]        ARSIZE_M2,
    input [`AXI_BURST_BITS-1:0]       ARBURST_M2,
    input                             ARVALID_M2,
    output logic                      ARREADY_M2,
    output logic [`AXI_ID_BITS-1:0]   RID_M2,
    output logic [`AXI_DATA_BITS-1:0] RDATA_M2,
    output logic [`AXI_RESP_BITS-1:0] RRESP_M2,
    output logic                      RLAST_M2,
    output logic                      RVALID_M2,
    input                             RREADY_M2,
    //SLAVE INTERFACE
    // S0
    // READ
    output logic [`AXI_IDS_BITS-1:0]  ARID_S0,
    output [`AXI_ADDR_BITS-1:0]       ARADDR_S0,
    output [`AXI_LEN_BITS-1:0]        ARLEN_S0,
    output [`AXI_SIZE_BITS-1:0]       ARSIZE_S0,
    output [`AXI_BURST_BITS-1:0]      ARBURST_S0,
    output logic                      ARVALID_S0,
    input                             ARREADY_S0,
    input [`AXI_IDS_BITS-1:0]         RID_S0,
    input [`AXI_DATA_BITS-1:0]        RDATA_S0,
    input [`AXI_RESP_BITS-1:0]        RRESP_S0,
    input                             RLAST_S0,
    input                             RVALID_S0,
    output logic                      RREADY_S0,
    // S1
    // WRITE
    output logic [`AXI_IDS_BITS-1:0]  AWID_S1,
    output [`AXI_ADDR_BITS-1:0]       AWADDR_S1,
    output [`AXI_LEN_BITS-1:0]        AWLEN_S1,
    output [`AXI_SIZE_BITS-1:0]       AWSIZE_S1,
    output [`AXI_BURST_BITS-1:0]      AWBURST_S1,
    output logic                      AWVALID_S1,
    input                             AWREADY_S1,
    output logic [`AXI_DATA_BITS-1:0] WDATA_S1,
    output logic [`AXI_STRB_BITS-1:0] WSTRB_S1,
    output logic                      WLAST_S1,
    output logic                      WVALID_S1,
    input                             WREADY_S1,
    input [`AXI_IDS_BITS-1:0]         BID_S1,
    input [`AXI_RESP_BITS-1:0]        BRESP_S1,
    input                             BVALID_S1,
    output logic                      BREADY_S1,
    // READ
    output logic [`AXI_IDS_BITS-1:0]  ARID_S1,
    output [`AXI_ADDR_BITS-1:0]       ARADDR_S1,
    output [`AXI_LEN_BITS-1:0]        ARLEN_S1,
    output [`AXI_SIZE_BITS-1:0]       ARSIZE_S1,
    output [`AXI_BURST_BITS-1:0]      ARBURST_S1,
    output logic                      ARVALID_S1,
    input                             ARREADY_S1,
    input [`AXI_IDS_BITS-1:0]         RID_S1,
    input [`AXI_DATA_BITS-1:0]        RDATA_S1,
    input [`AXI_RESP_BITS-1:0]        RRESP_S1,
    input                             RLAST_S1,
    input                             RVALID_S1,
    output logic                      RREADY_S1,
    // S2
    // WRITE
    output logic [`AXI_IDS_BITS-1:0]  AWID_S2,
    output [`AXI_ADDR_BITS-1:0]       AWADDR_S2,
    output [`AXI_LEN_BITS-1:0]        AWLEN_S2,
    output [`AXI_SIZE_BITS-1:0]       AWSIZE_S2,
    output [`AXI_BURST_BITS-1:0]      AWBURST_S2,
    output logic                      AWVALID_S2,
    input                             AWREADY_S2,
    output logic [`AXI_DATA_BITS-1:0] WDATA_S2,
    output logic [`AXI_STRB_BITS-1:0] WSTRB_S2,
    output logic                      WLAST_S2,
    output logic                      WVALID_S2,
    input                             WREADY_S2,
    input [`AXI_IDS_BITS-1:0]         BID_S2,
    input [`AXI_RESP_BITS-1:0]        BRESP_S2,
    input                             BVALID_S2,
    output logic                      BREADY_S2,
    // READ
    output logic [`AXI_IDS_BITS-1:0]  ARID_S2,
    output [`AXI_ADDR_BITS-1:0]       ARADDR_S2,
    output [`AXI_LEN_BITS-1:0]        ARLEN_S2,
    output [`AXI_SIZE_BITS-1:0]       ARSIZE_S2,
    output [`AXI_BURST_BITS-1:0]      ARBURST_S2,
    output logic                      ARVALID_S2,
    input                             ARREADY_S2,
    input [`AXI_IDS_BITS-1:0]         RID_S2,
    input [`AXI_DATA_BITS-1:0]        RDATA_S2,
    input [`AXI_RESP_BITS-1:0]        RRESP_S2,
    input                             RLAST_S2,
    input                             RVALID_S2,
    output logic                      RREADY_S2,
    // S3
    // WRITE
    output logic [`AXI_IDS_BITS-1:0]  AWID_S3,
    output [`AXI_ADDR_BITS-1:0]       AWADDR_S3,
    output [`AXI_LEN_BITS-1:0]        AWLEN_S3,
    output [`AXI_SIZE_BITS-1:0]       AWSIZE_S3,
    output [`AXI_BURST_BITS-1:0]      AWBURST_S3,
    output logic                      AWVALID_S3,
    input                             AWREADY_S3,
    output logic [`AXI_DATA_BITS-1:0] WDATA_S3,
    output logic [`AXI_STRB_BITS-1:0] WSTRB_S3,
    output logic                      WLAST_S3,
    output logic                      WVALID_S3,
    input                             WREADY_S3,
    input [`AXI_IDS_BITS-1:0]         BID_S3,
    input [`AXI_RESP_BITS-1:0]        BRESP_S3,
    input                             BVALID_S3,
    output  logic                     BREADY_S3,
    // READ
    output logic [`AXI_IDS_BITS-1:0]  ARID_S3,
    output [`AXI_ADDR_BITS-1:0]       ARADDR_S3,
    output [`AXI_LEN_BITS-1:0]        ARLEN_S3,
    output [`AXI_SIZE_BITS-1:0]       ARSIZE_S3,
    output [`AXI_BURST_BITS-1:0]      ARBURST_S3,
    output logic                      ARVALID_S3,
    input                             ARREADY_S3,
    input [`AXI_IDS_BITS-1:0]         RID_S3,
    input [`AXI_DATA_BITS-1:0]        RDATA_S3,
    input [`AXI_RESP_BITS-1:0]        RRESP_S3,
    input                             RLAST_S3,
    input                             RVALID_S3,
    output logic                      RREADY_S3,
    // S4
    // WRITE
    output logic [`AXI_IDS_BITS-1:0]  AWID_S4,
    output [`AXI_ADDR_BITS-1:0]       AWADDR_S4,
    output [`AXI_LEN_BITS-1:0]        AWLEN_S4,
    output [`AXI_SIZE_BITS-1:0]       AWSIZE_S4,
    output [`AXI_BURST_BITS-1:0]      AWBURST_S4,
    output logic                      AWVALID_S4,
    input                             AWREADY_S4,
    output logic [`AXI_DATA_BITS-1:0] WDATA_S4,
    output logic [`AXI_STRB_BITS-1:0] WSTRB_S4,
    output logic                      WLAST_S4,
    output logic                      WVALID_S4,
    input                             WREADY_S4,
    input [`AXI_IDS_BITS-1:0]         BID_S4,
    input [`AXI_RESP_BITS-1:0]        BRESP_S4,
    input                             BVALID_S4,
    output logic                      BREADY_S4,
    // READ
    output logic [`AXI_IDS_BITS-1:0]  ARID_S4,
    output [`AXI_ADDR_BITS-1:0]       ARADDR_S4,
    output [`AXI_LEN_BITS-1:0]        ARLEN_S4,
    output [`AXI_SIZE_BITS-1:0]       ARSIZE_S4,
    output [`AXI_BURST_BITS-1:0]      ARBURST_S4,
    output logic                      ARVALID_S4,
    input                             ARREADY_S4,
    input [`AXI_IDS_BITS-1:0]         RID_S4,
    input [`AXI_DATA_BITS-1:0]        RDATA_S4,
    input [`AXI_RESP_BITS-1:0]        RRESP_S4,
    input                             RLAST_S4,
    input                             RVALID_S4,
    output logic                      RREADY_S4,
    // S5
    // WRITE
    output logic [`AXI_IDS_BITS-1:0]  AWID_S5,
    output [`AXI_ADDR_BITS-1:0]       AWADDR_S5,
    output [`AXI_LEN_BITS-1:0]        AWLEN_S5,
    output [`AXI_SIZE_BITS-1:0]       AWSIZE_S5,
    output [`AXI_BURST_BITS-1:0]      AWBURST_S5,
    output logic                      AWVALID_S5,
    input                             AWREADY_S5,
    output logic [`AXI_DATA_BITS-1:0] WDATA_S5,
    output logic [`AXI_STRB_BITS-1:0] WSTRB_S5,
    output logic                      WLAST_S5,
    output logic                      WVALID_S5,
    input                             WREADY_S5,
    input [`AXI_IDS_BITS-1:0]         BID_S5,
    input [`AXI_RESP_BITS-1:0]        BRESP_S5,
    input                             BVALID_S5,
    output logic                      BREADY_S5,
    // READ
    output logic [`AXI_IDS_BITS-1:0]  ARID_S5,
    output [`AXI_ADDR_BITS-1:0]       ARADDR_S5,
    output [`AXI_LEN_BITS-1:0]        ARLEN_S5,
    output [`AXI_SIZE_BITS-1:0]       ARSIZE_S5,
    output [`AXI_BURST_BITS-1:0]      ARBURST_S5,
    output logic                      ARVALID_S5,
    input                             ARREADY_S5,
    input [`AXI_IDS_BITS-1:0]         RID_S5,
    input [`AXI_DATA_BITS-1:0]        RDATA_S5,
    input [`AXI_RESP_BITS-1:0]        RRESP_S5,
    input                             RLAST_S5,
    input                             RVALID_S5,
    output logic                      RREADY_S5,
    // S6
    // WRITE
    output logic [`AXI_IDS_BITS-1:0]  AWID_S6,
    output [`AXI_ADDR_BITS-1:0]       AWADDR_S6,
    output [`AXI_LEN_BITS-1:0]        AWLEN_S6,
    output [`AXI_SIZE_BITS-1:0]       AWSIZE_S6,
    output [`AXI_BURST_BITS-1:0]      AWBURST_S6,
    output logic                      AWVALID_S6,
    input                             AWREADY_S6,
    output logic [`AXI_DATA_BITS-1:0] WDATA_S6,
    output logic [`AXI_STRB_BITS-1:0] WSTRB_S6,
    output logic                      WLAST_S6,
    output logic                      WVALID_S6,
    input                             WREADY_S6,
    input [`AXI_IDS_BITS-1:0]         BID_S6,
    input [`AXI_RESP_BITS-1:0]        BRESP_S6,
    input                             BVALID_S6,
    output logic                      BREADY_S6,
    // READ
    output logic [`AXI_IDS_BITS-1:0]  ARID_S6,
    output [`AXI_ADDR_BITS-1:0]       ARADDR_S6,
    output [`AXI_LEN_BITS-1:0]        ARLEN_S6,
    output [`AXI_SIZE_BITS-1:0]       ARSIZE_S6,
    output [`AXI_BURST_BITS-1:0]      ARBURST_S6,
    output logic                      ARVALID_S6,
    input                             ARREADY_S6,
    input [`AXI_IDS_BITS-1:0]         RID_S6,
    input [`AXI_DATA_BITS-1:0]        RDATA_S6,
    input [`AXI_RESP_BITS-1:0]        RRESP_S6,
    input                             RLAST_S6,
    input                             RVALID_S6,
    output logic                      RREADY_S6,
    // S7
    // WRITE
    output logic [`AXI_IDS_BITS-1:0]  AWID_S7,
    output [`AXI_ADDR_BITS-1:0]       AWADDR_S7,
    output [`AXI_LEN_BITS-1:0]        AWLEN_S7,
    output [`AXI_SIZE_BITS-1:0]       AWSIZE_S7,
    output [`AXI_BURST_BITS-1:0]      AWBURST_S7,
    output logic                      AWVALID_S7,
    input                             AWREADY_S7,
    output logic [`AXI_DATA_BITS-1:0] WDATA_S7,
    output logic [`AXI_STRB_BITS-1:0] WSTRB_S7,
    output logic                      WLAST_S7,
    output logic                      WVALID_S7,
    input                             WREADY_S7,
    input [`AXI_IDS_BITS-1:0]         BID_S7,
    input [`AXI_RESP_BITS-1:0]        BRESP_S7,
    input                             BVALID_S7,
    output logic                      BREADY_S7,
    // READ
    output logic [`AXI_IDS_BITS-1:0]  ARID_S7,
    output [`AXI_ADDR_BITS-1:0]       ARADDR_S7,
    output [`AXI_LEN_BITS-1:0]        ARLEN_S7,
    output [`AXI_SIZE_BITS-1:0]       ARSIZE_S7,
    output [`AXI_BURST_BITS-1:0]      ARBURST_S7,
    output logic                      ARVALID_S7,
    input                             ARREADY_S7,
    input [`AXI_IDS_BITS-1:0]         RID_S7,
    input [`AXI_DATA_BITS-1:0]        RDATA_S7,
    input [`AXI_RESP_BITS-1:0]        RRESP_S7,
    input                             RLAST_S7,
    input                             RVALID_S7,
    output logic                      RREADY_S7
);

// ROM      0x0000_0000 ~ 0x0000_1FFF
// IM       0x0001_0000 ~ 0x0001_FFFF
// DM       0x0002_0000 ~ 0x0002_FFFF
// Sctrl    0x1000_0000 ~ 0x1000_03FF
// DRAM     0x2000_0000 ~ 0x201F_FFFF
// DMA      0x3000_0000 ~ 0x3000_0FFF
// TPU      0x3000_1000 ~ 0x3000_100F

AXI_rd AXI_rd0(
    .ACLK(ACLK),
    .ARESETn(ARESETn),
    //SLAVE INTERFACE FOR MASTERS
    // M0
    .ARID_M0(ARID_M0),
    .ARADDR_M0(ARADDR_M0),
    .ARLEN_M0(ARLEN_M0),
    .ARSIZE_M0(ARSIZE_M0),
    .ARBURST_M0(ARBURST_M0),
    .ARVALID_M0(ARVALID_M0),
    .ARREADY_M0(ARREADY_M0),
    .RID_M0(RID_M0),
    .RDATA_M0(RDATA_M0),
    .RRESP_M0(RRESP_M0),
    .RLAST_M0(RLAST_M0),
    .RVALID_M0(RVALID_M0),
    .RREADY_M0(RREADY_M0),
    
    // M1
    .ARID_M1(ARID_M1),
    .ARADDR_M1(ARADDR_M1),
    .ARLEN_M1(ARLEN_M1),
    .ARSIZE_M1(ARSIZE_M1),
    .ARBURST_M1(ARBURST_M1),
    .ARVALID_M1(ARVALID_M1),
    .ARREADY_M1(ARREADY_M1),
    .RID_M1(RID_M1),
    .RDATA_M1(RDATA_M1),
    .RRESP_M1(RRESP_M1),
    .RLAST_M1(RLAST_M1),
    .RVALID_M1(RVALID_M1),
    .RREADY_M1(RREADY_M1),

    // M2
    .ARID_M2(ARID_M2),
    .ARADDR_M2(ARADDR_M2),
    .ARLEN_M2(ARLEN_M2),
    .ARSIZE_M2(ARSIZE_M2),
    .ARBURST_M2(ARBURST_M2),
    .ARVALID_M2(ARVALID_M2),
    .ARREADY_M2(ARREADY_M2),
    .RID_M2(RID_M2),
    .RDATA_M2(RDATA_M2),
    .RRESP_M2(RRESP_M2),
    .RLAST_M2(RLAST_M2),
    .RVALID_M2(RVALID_M2),
    .RREADY_M2(RREADY_M2),

    //MASTER INTERFACE FOR SLAVES
    // S0
    .ARID_S0(ARID_S0),
    .ARADDR_S0(ARADDR_S0),
    .ARLEN_S0(ARLEN_S0),
    .ARSIZE_S0(ARSIZE_S0),
    .ARBURST_S0(ARBURST_S0),
    .ARVALID_S0(ARVALID_S0),
    .ARREADY_S0(ARREADY_S0),
    .RID_S0(RID_S0),
    .RDATA_S0(RDATA_S0),
    .RRESP_S0(RRESP_S0),
    .RLAST_S0(RLAST_S0),
    .RVALID_S0(RVALID_S0),
    .RREADY_S0(RREADY_S0),

    // S1
    .ARID_S1(ARID_S1),
    .ARADDR_S1(ARADDR_S1),
    .ARLEN_S1(ARLEN_S1),
    .ARSIZE_S1(ARSIZE_S1),
    .ARBURST_S1(ARBURST_S1),
    .ARVALID_S1(ARVALID_S1),
    .ARREADY_S1(ARREADY_S1),
    .RID_S1(RID_S1),
    .RDATA_S1(RDATA_S1),
    .RRESP_S1(RRESP_S1),
    .RLAST_S1(RLAST_S1),
    .RVALID_S1(RVALID_S1),
    .RREADY_S1(RREADY_S1),

    // S2
    .ARID_S2(ARID_S2),
    .ARADDR_S2(ARADDR_S2),
    .ARLEN_S2(ARLEN_S2),
    .ARSIZE_S2(ARSIZE_S2),
    .ARBURST_S2(ARBURST_S2),
    .ARVALID_S2(ARVALID_S2),
    .ARREADY_S2(ARREADY_S2),
    .RID_S2(RID_S2),
    .RDATA_S2(RDATA_S2),
    .RRESP_S2(RRESP_S2),
    .RLAST_S2(RLAST_S2),
    .RVALID_S2(RVALID_S2),
    .RREADY_S2(RREADY_S2),

    // S3
    .ARID_S3(ARID_S3),
    .ARADDR_S3(ARADDR_S3),
    .ARLEN_S3(ARLEN_S3),
    .ARSIZE_S3(ARSIZE_S3),
    .ARBURST_S3(ARBURST_S3),
    .ARVALID_S3(ARVALID_S3),
    .ARREADY_S3(ARREADY_S3),
    .RID_S3(RID_S3),
    .RDATA_S3(RDATA_S3),
    .RRESP_S3(RRESP_S3),
    .RLAST_S3(RLAST_S3),
    .RVALID_S3(RVALID_S3),
    .RREADY_S3(RREADY_S3),

    // S4
    .ARID_S4(ARID_S4),
    .ARADDR_S4(ARADDR_S4),
    .ARLEN_S4(ARLEN_S4),
    .ARSIZE_S4(ARSIZE_S4),
    .ARBURST_S4(ARBURST_S4),
    .ARVALID_S4(ARVALID_S4),
    .ARREADY_S4(ARREADY_S4),
    .RID_S4(RID_S4),
    .RDATA_S4(RDATA_S4),
    .RRESP_S4(RRESP_S4),
    .RLAST_S4(RLAST_S4),
    .RVALID_S4(RVALID_S4),
    .RREADY_S4(RREADY_S4),

    // S5
    .ARID_S5(ARID_S5),
    .ARADDR_S5(ARADDR_S5),
    .ARLEN_S5(ARLEN_S5),
    .ARSIZE_S5(ARSIZE_S5),
    .ARBURST_S5(ARBURST_S5),
    .ARVALID_S5(ARVALID_S5),
    .ARREADY_S5(ARREADY_S5),
    .RID_S5(RID_S5),
    .RDATA_S5(RDATA_S5),
    .RRESP_S5(RRESP_S5),
    .RLAST_S5(RLAST_S5),
    .RVALID_S5(RVALID_S5),
    .RREADY_S5(RREADY_S5),

    // S6
    .ARID_S6(ARID_S6),
    .ARADDR_S6(ARADDR_S6),
    .ARLEN_S6(ARLEN_S6),
    .ARSIZE_S6(ARSIZE_S6),
    .ARBURST_S6(ARBURST_S6),
    .ARVALID_S6(ARVALID_S6),
    .ARREADY_S6(ARREADY_S6),
    .RID_S6(RID_S6),
    .RDATA_S6(RDATA_S6),
    .RRESP_S6(RRESP_S6),
    .RLAST_S6(RLAST_S6),
    .RVALID_S6(RVALID_S6),
    .RREADY_S6(RREADY_S6),

    // S7
    .ARID_S7(ARID_S7),
    .ARADDR_S7(ARADDR_S7),
    .ARLEN_S7(ARLEN_S7),
    .ARSIZE_S7(ARSIZE_S7),
    .ARBURST_S7(ARBURST_S7),
    .ARVALID_S7(ARVALID_S7),
    .ARREADY_S7(ARREADY_S7),
    .RID_S7(RID_S7),
    .RDATA_S7(RDATA_S7),
    .RRESP_S7(RRESP_S7),
    .RLAST_S7(RLAST_S7),
    .RVALID_S7(RVALID_S7),
    .RREADY_S7(RREADY_S7)
);

AXI_wr AXI_wr0(
    .ACLK(ACLK),
    .ARESETn(ARESETn),

    //SLAVE INTERFACE FOR MASTERS
    // M1
    .AWID_M1(AWID_M1),
    .AWADDR_M1(AWADDR_M1),
    .AWLEN_M1(AWLEN_M1),
    .AWSIZE_M1(AWSIZE_M1),
    .AWBURST_M1(AWBURST_M1),
    .AWVALID_M1(AWVALID_M1),
    .AWREADY_M1(AWREADY_M1),
    .WDATA_M1(WDATA_M1),
    .WSTRB_M1(WSTRB_M1),
    .WLAST_M1(WLAST_M1),
    .WVALID_M1(WVALID_M1),
    .WREADY_M1(WREADY_M1),
    .BID_M1(BID_M1),
    .BRESP_M1(BRESP_M1),
    .BVALID_M1(BVALID_M1),
    .BREADY_M1(BREADY_M1),

    // M2
    .AWID_M2(AWID_M2),
    .AWADDR_M2(AWADDR_M2),
    .AWLEN_M2(AWLEN_M2),
    .AWSIZE_M2(AWSIZE_M2),
    .AWBURST_M2(AWBURST_M2),
    .AWVALID_M2(AWVALID_M2),
    .AWREADY_M2(AWREADY_M2),
    .WDATA_M2(WDATA_M2),
    .WSTRB_M2(WSTRB_M2),
    .WLAST_M2(WLAST_M2),
    .WVALID_M2(WVALID_M2),
    .WREADY_M2(WREADY_M2),
    .BID_M2(BID_M2),
    .BRESP_M2(BRESP_M2),
    .BVALID_M2(BVALID_M2),
    .BREADY_M2(BREADY_M2),

    //MASTER INTERFACE FOR SLAVES
    // S1
    .AWID_S1(AWID_S1),
    .AWADDR_S1(AWADDR_S1),
    .AWLEN_S1(AWLEN_S1),
    .AWSIZE_S1(AWSIZE_S1),
    .AWBURST_S1(AWBURST_S1),
    .AWVALID_S1(AWVALID_S1),
    .AWREADY_S1(AWREADY_S1),
    .WDATA_S1(WDATA_S1),
    .WSTRB_S1(WSTRB_S1),
    .WLAST_S1(WLAST_S1),
    .WVALID_S1(WVALID_S1),
    .WREADY_S1(WREADY_S1),
    .BID_S1(BID_S1),
    .BRESP_S1(BRESP_S1),
    .BVALID_S1(BVALID_S1),
    .BREADY_S1(BREADY_S1),

    // S2
    .AWID_S2(AWID_S2),
    .AWADDR_S2(AWADDR_S2),
    .AWLEN_S2(AWLEN_S2),
    .AWSIZE_S2(AWSIZE_S2),
    .AWBURST_S2(AWBURST_S2),
    .AWVALID_S2(AWVALID_S2),
    .AWREADY_S2(AWREADY_S2),
    .WDATA_S2(WDATA_S2),
    .WSTRB_S2(WSTRB_S2),
    .WLAST_S2(WLAST_S2),
    .WVALID_S2(WVALID_S2),
    .WREADY_S2(WREADY_S2),
    .BID_S2(BID_S2),
    .BRESP_S2(BRESP_S2),
    .BVALID_S2(BVALID_S2),
    .BREADY_S2(BREADY_S2),

    // S3
    .AWID_S3(AWID_S3),
    .AWADDR_S3(AWADDR_S3),
    .AWLEN_S3(AWLEN_S3),
    .AWSIZE_S3(AWSIZE_S3),
    .AWBURST_S3(AWBURST_S3),
    .AWVALID_S3(AWVALID_S3),
    .AWREADY_S3(AWREADY_S3),
    .WDATA_S3(WDATA_S3),
    .WSTRB_S3(WSTRB_S3),
    .WLAST_S3(WLAST_S3),
    .WVALID_S3(WVALID_S3),
    .WREADY_S3(WREADY_S3),
    .BID_S3(BID_S3),
    .BRESP_S3(BRESP_S3),
    .BVALID_S3(BVALID_S3),
    .BREADY_S3(BREADY_S3),

    // S4
    .AWID_S4(AWID_S4),
    .AWADDR_S4(AWADDR_S4),
    .AWLEN_S4(AWLEN_S4),
    .AWSIZE_S4(AWSIZE_S4),
    .AWBURST_S4(AWBURST_S4),
    .AWVALID_S4(AWVALID_S4),
    .AWREADY_S4(AWREADY_S4),
    .WDATA_S4(WDATA_S4),
    .WSTRB_S4(WSTRB_S4),
    .WLAST_S4(WLAST_S4),
    .WVALID_S4(WVALID_S4),
    .WREADY_S4(WREADY_S4),
    .BID_S4(BID_S4),
    .BRESP_S4(BRESP_S4),
    .BVALID_S4(BVALID_S4),
    .BREADY_S4(BREADY_S4),

    // S5
    .AWID_S5(AWID_S5),
    .AWADDR_S5(AWADDR_S5),
    .AWLEN_S5(AWLEN_S5),
    .AWSIZE_S5(AWSIZE_S5),
    .AWBURST_S5(AWBURST_S5),
    .AWVALID_S5(AWVALID_S5),
    .AWREADY_S5(AWREADY_S5),
    .WDATA_S5(WDATA_S5),
    .WSTRB_S5(WSTRB_S5),
    .WLAST_S5(WLAST_S5),
    .WVALID_S5(WVALID_S5),
    .WREADY_S5(WREADY_S5),
    .BID_S5(BID_S5),
    .BRESP_S5(BRESP_S5),
    .BVALID_S5(BVALID_S5),
    .BREADY_S5(BREADY_S5),

    // S6
    .AWID_S6(AWID_S6),
    .AWADDR_S6(AWADDR_S6),
    .AWLEN_S6(AWLEN_S6),
    .AWSIZE_S6(AWSIZE_S6),
    .AWBURST_S6(AWBURST_S6),
    .AWVALID_S6(AWVALID_S6),
    .AWREADY_S6(AWREADY_S6),
    .WDATA_S6(WDATA_S6),
    .WSTRB_S6(WSTRB_S6),
    .WLAST_S6(WLAST_S6),
    .WVALID_S6(WVALID_S6),
    .WREADY_S6(WREADY_S6),
    .BID_S6(BID_S6),
    .BRESP_S6(BRESP_S6),
    .BVALID_S6(BVALID_S6),
    .BREADY_S6(BREADY_S6),

    // S7
    .AWID_S7(AWID_S7),
    .AWADDR_S7(AWADDR_S7),
    .AWLEN_S7(AWLEN_S7),
    .AWSIZE_S7(AWSIZE_S7),
    .AWBURST_S7(AWBURST_S7),
    .AWVALID_S7(AWVALID_S7),
    .AWREADY_S7(AWREADY_S7),
    .WDATA_S7(WDATA_S7),
    .WSTRB_S7(WSTRB_S7),
    .WLAST_S7(WLAST_S7),
    .WVALID_S7(WVALID_S7),
    .WREADY_S7(WREADY_S7),
    .BID_S7(BID_S7),
    .BRESP_S7(BRESP_S7),
    .BVALID_S7(BVALID_S7),
    .BREADY_S7(BREADY_S7)
);


endmodule
